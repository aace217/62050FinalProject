`timescale 1ns / 1ps
`default_nettype none

module note_storing_pixel_addressing(
    input wire rst_in,
    input wire clk_in,
);



endmodule
`default_nettype wire
