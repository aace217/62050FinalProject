`timescale 1ns / 1ps
`default_nettype none
module midi_decode(
    input wire midi_Data_in,
    input wire rst_in,
    input wire clk_in,
    output logic [34:0] velocity,
    output logic [34:0] received_note

);
    // calculate 
endmodule
`default_nettype wire
