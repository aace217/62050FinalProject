`timescale 1ns / 1ps
`default_nettype none

module baton_tracker(
    input wire [10:0] x_com_in,
    input wire [9:0] y_com_in,
    input wire measure_in,
    input wire rst_in,
    input wire clk_camera_in,
    output logic change_out
)
endmodule
`default_nettype wire
